module adder#(
    parameter DATA_WIDTH = 32,
    parameter ADDRESS_SIZE = 8
)
(
    input ACLK  // Global clock signal
    input ARESETn //Global reset signal, of type active LOW 
);

endmodule